module tb_comb_Y2;
    wire Y;
    reg A,B,C,D;

    comb_Y2 a(Y, A, B, C, D);

integer k;

    initial 
    begin
        for ( k=1; k<16; k=k+1 )
        begin
            {A,B,C,D} = k;
            #5;
        end
    end

    initial
        $monitor("At time %4t, A=%b, B=%b, C=%b, D=%b, Y=%b",
                    $time, A, B, C, D, Y);
endmodule
