module tb_shift_counter;
    wire [7:0] count;
    reg clk,reset;

    shift_counter a(count,clk,reset);

    initial
    begin
        reset = 1'b0;
        #50 reset = 1'b1;
        #15 reset = 1'b0; 
    end

    initial
    begin
        clk = 1'b0;
        forever #5 clk = ~clk;
    end

    initial
        $monitor("At time %4t, reset=%b, count=%b",
                    $time, reset, count);
endmodule
